library ieee;
use ieee.std_logic_1164.all;


entity elevator_sim is
  port(

      );


end elevator_sim;
